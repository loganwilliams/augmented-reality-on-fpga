// Logan Williams


module pt_fetcher(
		  // STANDARD INPUTS
		  input 	    clock,
		  input 	    reset,
		  // TO AND FROM PROJECTIVE_TRANSFORM
		  input 	    pt_flag,
		  input [9:0] 	    pt_x,
		  input [8:0] 	    pt_y,
		  input [17:0] 	    pt_pixel,
		  output 	    done_pt,
		  // TO AND FROM MEMORY_INTERFACE
		  input [35:0] 	    ptf_pixel_read,
		  input 	    done_ptf,
		  output reg [9:0]  ptf_x,
		  output reg [8:0]  ptf_y,
		  output reg 	    ptf_flag,
		  output reg 	    ptf_wr,
		  output reg [35:0] ptf_pixel_write);
   

   reg [17:0] 			    pt_pixel_buffer [0:1];
   reg [9:0] 			    pt_pixel_x [0:1];
   reg [8:0] 			    pt_pixel_y [0:1];
   reg 				    haspixel;
   reg [1:0] 			    state;
   

   assign done_pt = done_ptf & (~state[1]);

   always @(posedge clock) begin
      if (reset) begin
	 // reset everything to its initial state
	 state <= 2'b00;
	 pt_pixel_buffer[0] <= 0;
	 pt_pixel_buffer[1] <= 0;
	 pt_pixel_x[0] <= 0;
	 pt_pixel_x[1] <= 0;
	 pt_pixel_y[0] <= 0;
	 pt_pixel_y[1] <= 0;
	 haspixel <= 0;
	 
      end
      
      case (state)
	2'b00: begin
	   if (pt_flag) begin
	      pt_pixel_buffer[0] <= pt_pixel;
	      pt_pixel_x[0] <= pt_x;
	      pt_pixel_y[0] <= pt_y;
	      haspixel = 1;
	   end

	   if (done_ptf & haspixel) begin
	      ptf_x <= pt_x;
	      ptf_y <= pt_y;
	      ptf_wr <= 0;
	      ptf_flag <= 1;
	      state <= 2'b01;
	      haspixel <= 0;
	      
	   end 
	end

	2'b01: begin
	   if (pt_flag) begin
	      pt_pixel_buffer[1] <= pt_pixel;
	      pt_pixel_x[1] <= pt_x;
	      pt_pixel_y[1] <= pt_y;
	      haspixel = 1;
	      
	   end

	   if (done_ptf & haspixel) begin
	      ptf_x <= pt_x;
	      ptf_y <= pt_y;
	      ptf_wr <= 0;
	      ptf_flag <= 1;
	      state <= 2'b10;
	      haspixel <= 0;
	   end 
	end

	2'b10: begin

	   
	   // catch the case where both pixels are in the same address
	   if ((pt_pixel_x[0] >> 1) == (pt_pixel_x[1] >> 1) & 
	       (pt_pixel_y[0] == pt_pixel_y[1]) & (pt_pixel_x[0] != pt_pixel_x[1])) begin
	      if (pt_pixel_x[0] < pt_pixel_x[1]) begin
		 ptf_pixel_write <= {pt_pixel_buffer[1],pt_pixel_buffer[0]};
		 ptf_x <= pt_pixel_x[0];
		 ptf_y <= pt_pixel_y[0];
	      end else begin
		 ptf_pixel_write <= {pt_pixel_buffer[0],pt_pixel_buffer[1]};
		 ptf_x <= pt_pixel_x[1];
		 ptf_y <= pt_pixel_y[1];
	      end

	      // skip the fourth state
	      state <= 2'b00;
	      ptf_flag <= 1;
	      ptf_wr <= 1;
	      
	   end else begin // if ((pt_pixel_x[0] >> 1) == (pt_pixel_x[1] >> 1) &...
	      
	      
	      // concatenate normally
	      if (pt_pixel_x[0][0]) ptf_pixel_write <= {ptf_pixel_read[35:18], pt_pixel_buffer[0]};
	      else ptf_pixel_write <= {pt_pixel_buffer[0], ptf_pixel_read[17:0]};
	      
	      
	      // send write for new pixel pair
	      ptf_x <= pt_pixel_x[0];
	      ptf_y <= pt_pixel_y[0];
	      ptf_flag <= 1;
	      ptf_wr <= 1;
	      
	      // go to next state
	      state <= 2'b11;
	   end
	end

	2'b11: begin
	   // concatenate

	   if (pt_pixel_x[1][0]) ptf_pixel_write <= {ptf_pixel_read[35:18], pt_pixel_buffer[1]};
	   else ptf_pixel_write <= {pt_pixel_buffer[1], ptf_pixel_read[17:0]};

	   // send write for new pixel pair

	   ptf_x <= pt_pixel_x[1];
	   ptf_y <= pt_pixel_y[1];
	   ptf_flag <= 1;
	   ptf_wr <= 1;

	   state <= 2'b00;
	   
	end
      endcase // case state
   end // always @ (posedge clock)
   
endmodule // pt_fetcher