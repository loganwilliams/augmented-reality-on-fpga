library verilog;
use verilog.vl_types.all;
entity test_pt_fetcher is
end test_pt_fetcher;
