library verilog;
use verilog.vl_types.all;
entity test_ntsc_clean is
end test_ntsc_clean;
