library verilog;
use verilog.vl_types.all;
entity projective_transform_test is
end projective_transform_test;
